library verilog;
use verilog.vl_types.all;
entity \testbench__lhlb\ is
end \testbench__lhlb\;
