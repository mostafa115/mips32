library verilog;
use verilog.vl_types.all;
entity \testbench__andi\ is
end \testbench__andi\;
