library verilog;
use verilog.vl_types.all;
entity testbench_lbu is
end testbench_lbu;
